// Automatically synthesized high-speed adder (AHSA) of size 32-bits

module ahsa_32b ( a, b, sum );
  input [31:0] a;
  input [31:0] b;
  output [32:0] sum;
  wire   \intadd_0/n38 , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314;
  assign sum[32] = \intadd_0/n38 ;

  NOR2X0_HVT U35 ( .A1(a[21]), .A2(b[21]), .Y(n153) );
  NOR2X0_HVT U36 ( .A1(a[20]), .A2(b[20]), .Y(n147) );
  NOR2X0_HVT U37 ( .A1(n153), .A2(n147), .Y(n139) );
  NOR2X0_HVT U38 ( .A1(a[23]), .A2(b[23]), .Y(n133) );
  NOR2X0_HVT U39 ( .A1(a[22]), .A2(b[22]), .Y(n142) );
  NOR2X0_HVT U40 ( .A1(n133), .A2(n142), .Y(n50) );
  NAND2X0_HVT U41 ( .A1(n139), .A2(n50), .Y(n52) );
  NOR2X0_HVT U42 ( .A1(a[17]), .A2(b[17]), .Y(n181) );
  NOR2X0_HVT U43 ( .A1(a[16]), .A2(b[16]), .Y(n186) );
  NOR2X0_HVT U44 ( .A1(n181), .A2(n186), .Y(n173) );
  NOR2X0_HVT U45 ( .A1(a[19]), .A2(b[19]), .Y(n168) );
  NOR2X0_HVT U46 ( .A1(a[18]), .A2(b[18]), .Y(n164) );
  NOR2X0_HVT U47 ( .A1(n168), .A2(n164), .Y(n48) );
  NAND2X0_HVT U48 ( .A1(n173), .A2(n48), .Y(n159) );
  NOR2X0_HVT U49 ( .A1(n52), .A2(n159), .Y(n193) );
  NOR2X0_HVT U50 ( .A1(b[29]), .A2(a[29]), .Y(n78) );
  NOR2X0_HVT U51 ( .A1(b[28]), .A2(a[28]), .Y(n87) );
  NOR2X0_HVT U52 ( .A1(n78), .A2(n87), .Y(n191) );
  NOR2X0_HVT U53 ( .A1(b[30]), .A2(a[30]), .Y(n190) );
  INVX1_HVT U54 ( .A(n190), .Y(n71) );
  NAND2X0_HVT U55 ( .A1(n191), .A2(n71), .Y(n57) );
  NOR2X0_HVT U56 ( .A1(a[25]), .A2(b[25]), .Y(n116) );
  NOR2X0_HVT U57 ( .A1(a[24]), .A2(b[24]), .Y(n112) );
  NOR2X0_HVT U58 ( .A1(n116), .A2(n112), .Y(n104) );
  NOR2X0_HVT U59 ( .A1(a[27]), .A2(b[27]), .Y(n98) );
  NOR2X0_HVT U60 ( .A1(a[26]), .A2(b[26]), .Y(n107) );
  NOR2X0_HVT U61 ( .A1(n98), .A2(n107), .Y(n54) );
  NAND2X0_HVT U62 ( .A1(n104), .A2(n54), .Y(n192) );
  NOR2X0_HVT U63 ( .A1(n57), .A2(n192), .Y(n59) );
  NAND2X0_HVT U64 ( .A1(n193), .A2(n59), .Y(n61) );
  NOR2X0_HVT U65 ( .A1(b[5]), .A2(a[5]), .Y(n289) );
  NOR2X0_HVT U66 ( .A1(b[4]), .A2(a[4]), .Y(n287) );
  NOR2X0_HVT U67 ( .A1(n289), .A2(n287), .Y(n276) );
  NOR2X0_HVT U68 ( .A1(b[7]), .A2(a[7]), .Y(n277) );
  NOR2X0_HVT U69 ( .A1(b[6]), .A2(a[6]), .Y(n282) );
  NOR2X0_HVT U70 ( .A1(n277), .A2(n282), .Y(n36) );
  NAND2X0_HVT U71 ( .A1(n276), .A2(n36), .Y(n38) );
  NAND2X0_HVT U72 ( .A1(a[0]), .A2(b[0]), .Y(n314) );
  NOR2X0_HVT U73 ( .A1(b[1]), .A2(a[1]), .Y(n309) );
  NAND2X0_HVT U74 ( .A1(a[1]), .A2(b[1]), .Y(n310) );
  OAI21X1_HVT U75 ( .A1(n314), .A2(n309), .A3(n310), .Y(n298) );
  NOR2X0_HVT U76 ( .A1(b[3]), .A2(a[3]), .Y(n299) );
  NOR2X0_HVT U77 ( .A1(b[2]), .A2(a[2]), .Y(n304) );
  NOR2X0_HVT U78 ( .A1(n299), .A2(n304), .Y(n34) );
  NAND2X0_HVT U79 ( .A1(a[2]), .A2(b[2]), .Y(n305) );
  NAND2X0_HVT U80 ( .A1(a[3]), .A2(b[3]), .Y(n300) );
  OAI21X1_HVT U81 ( .A1(n305), .A2(n299), .A3(n300), .Y(n33) );
  AOI21X1_HVT U82 ( .A1(n298), .A2(n34), .A3(n33), .Y(n274) );
  NAND2X0_HVT U83 ( .A1(a[4]), .A2(b[4]), .Y(n294) );
  NAND2X0_HVT U84 ( .A1(a[5]), .A2(b[5]), .Y(n290) );
  OAI21X1_HVT U85 ( .A1(n294), .A2(n289), .A3(n290), .Y(n275) );
  NAND2X0_HVT U86 ( .A1(a[6]), .A2(b[6]), .Y(n283) );
  NAND2X0_HVT U87 ( .A1(a[7]), .A2(b[7]), .Y(n278) );
  OAI21X1_HVT U88 ( .A1(n283), .A2(n277), .A3(n278), .Y(n35) );
  AOI21X1_HVT U89 ( .A1(n275), .A2(n36), .A3(n35), .Y(n37) );
  OAI21X1_HVT U90 ( .A1(n38), .A2(n274), .A3(n37), .Y(n210) );
  NOR2X0_HVT U91 ( .A1(a[13]), .A2(b[13]), .Y(n236) );
  NOR2X0_HVT U92 ( .A1(a[12]), .A2(b[12]), .Y(n230) );
  NOR2X0_HVT U93 ( .A1(n236), .A2(n230), .Y(n222) );
  NOR2X0_HVT U94 ( .A1(a[15]), .A2(b[15]), .Y(n216) );
  NOR2X0_HVT U95 ( .A1(a[14]), .A2(b[14]), .Y(n225) );
  NOR2X0_HVT U96 ( .A1(n216), .A2(n225), .Y(n42) );
  NAND2X0_HVT U97 ( .A1(n222), .A2(n42), .Y(n44) );
  NOR2X0_HVT U98 ( .A1(a[9]), .A2(b[9]), .Y(n264) );
  NOR2X0_HVT U99 ( .A1(a[8]), .A2(b[8]), .Y(n269) );
  NOR2X0_HVT U100 ( .A1(n264), .A2(n269), .Y(n256) );
  NOR2X0_HVT U101 ( .A1(a[11]), .A2(b[11]), .Y(n251) );
  NOR2X0_HVT U102 ( .A1(a[10]), .A2(b[10]), .Y(n247) );
  NOR2X0_HVT U103 ( .A1(n251), .A2(n247), .Y(n40) );
  NAND2X0_HVT U104 ( .A1(n256), .A2(n40), .Y(n242) );
  NOR2X0_HVT U105 ( .A1(n44), .A2(n242), .Y(n46) );
  NAND2X0_HVT U106 ( .A1(b[8]), .A2(a[8]), .Y(n270) );
  NAND2X0_HVT U107 ( .A1(b[9]), .A2(a[9]), .Y(n265) );
  OAI21X1_HVT U108 ( .A1(n270), .A2(n264), .A3(n265), .Y(n257) );
  NAND2X0_HVT U109 ( .A1(b[10]), .A2(a[10]), .Y(n260) );
  NAND2X0_HVT U110 ( .A1(b[11]), .A2(a[11]), .Y(n252) );
  OAI21X1_HVT U111 ( .A1(n260), .A2(n251), .A3(n252), .Y(n39) );
  AOI21X1_HVT U112 ( .A1(n257), .A2(n40), .A3(n39), .Y(n241) );
  NAND2X0_HVT U113 ( .A1(b[12]), .A2(a[12]), .Y(n243) );
  NAND2X0_HVT U114 ( .A1(b[13]), .A2(a[13]), .Y(n237) );
  OAI21X1_HVT U115 ( .A1(n243), .A2(n236), .A3(n237), .Y(n221) );
  NAND2X0_HVT U116 ( .A1(b[14]), .A2(a[14]), .Y(n226) );
  NAND2X0_HVT U117 ( .A1(b[15]), .A2(a[15]), .Y(n217) );
  OAI21X1_HVT U118 ( .A1(n226), .A2(n216), .A3(n217), .Y(n41) );
  AOI21X1_HVT U119 ( .A1(n221), .A2(n42), .A3(n41), .Y(n43) );
  OAI21X1_HVT U120 ( .A1(n44), .A2(n241), .A3(n43), .Y(n45) );
  AOI21X1_HVT U121 ( .A1(n210), .A2(n46), .A3(n45), .Y(n207) );
  NAND2X0_HVT U122 ( .A1(b[16]), .A2(a[16]), .Y(n187) );
  NAND2X0_HVT U123 ( .A1(b[17]), .A2(a[17]), .Y(n182) );
  OAI21X1_HVT U124 ( .A1(n187), .A2(n181), .A3(n182), .Y(n174) );
  NAND2X0_HVT U125 ( .A1(b[18]), .A2(a[18]), .Y(n177) );
  NAND2X0_HVT U126 ( .A1(b[19]), .A2(a[19]), .Y(n169) );
  OAI21X1_HVT U127 ( .A1(n177), .A2(n168), .A3(n169), .Y(n47) );
  AOI21X1_HVT U128 ( .A1(n174), .A2(n48), .A3(n47), .Y(n158) );
  NAND2X0_HVT U129 ( .A1(b[20]), .A2(a[20]), .Y(n160) );
  NAND2X0_HVT U130 ( .A1(b[21]), .A2(a[21]), .Y(n154) );
  OAI21X1_HVT U131 ( .A1(n160), .A2(n153), .A3(n154), .Y(n138) );
  NAND2X0_HVT U132 ( .A1(b[22]), .A2(a[22]), .Y(n143) );
  NAND2X0_HVT U133 ( .A1(b[23]), .A2(a[23]), .Y(n134) );
  OAI21X1_HVT U134 ( .A1(n143), .A2(n133), .A3(n134), .Y(n49) );
  AOI21X1_HVT U135 ( .A1(n138), .A2(n50), .A3(n49), .Y(n51) );
  OAI21X1_HVT U136 ( .A1(n52), .A2(n158), .A3(n51), .Y(n205) );
  NAND2X0_HVT U137 ( .A1(b[24]), .A2(a[24]), .Y(n123) );
  NAND2X0_HVT U138 ( .A1(b[25]), .A2(a[25]), .Y(n117) );
  OAI21X1_HVT U139 ( .A1(n123), .A2(n116), .A3(n117), .Y(n103) );
  NAND2X0_HVT U140 ( .A1(b[26]), .A2(a[26]), .Y(n108) );
  NAND2X0_HVT U141 ( .A1(b[27]), .A2(a[27]), .Y(n99) );
  OAI21X1_HVT U142 ( .A1(n108), .A2(n98), .A3(n99), .Y(n53) );
  AOI21X1_HVT U143 ( .A1(n103), .A2(n54), .A3(n53), .Y(n201) );
  NAND2X0_HVT U144 ( .A1(a[28]), .A2(b[28]), .Y(n88) );
  NAND2X0_HVT U145 ( .A1(a[29]), .A2(b[29]), .Y(n79) );
  OAI21X1_HVT U146 ( .A1(n88), .A2(n78), .A3(n79), .Y(n199) );
  NAND2X0_HVT U147 ( .A1(a[30]), .A2(b[30]), .Y(n196) );
  INVX1_HVT U148 ( .A(n196), .Y(n55) );
  AOI21X1_HVT U149 ( .A1(n199), .A2(n71), .A3(n55), .Y(n56) );
  OAI21X1_HVT U150 ( .A1(n57), .A2(n201), .A3(n56), .Y(n58) );
  AOI21X1_HVT U151 ( .A1(n205), .A2(n59), .A3(n58), .Y(n60) );
  OAI21X1_HVT U152 ( .A1(n61), .A2(n207), .A3(n60), .Y(n64) );
  NOR2X0_HVT U153 ( .A1(b[31]), .A2(a[31]), .Y(n195) );
  INVX1_HVT U154 ( .A(n195), .Y(n62) );
  NAND2X0_HVT U155 ( .A1(a[31]), .A2(b[31]), .Y(n194) );
  NAND2X0_HVT U156 ( .A1(n62), .A2(n194), .Y(n63) );
  XNOR2X1_HVT U157 ( .A1(n64), .A2(n63), .Y(sum[31]) );
  INVX1_HVT U158 ( .A(n191), .Y(n66) );
  NOR2X0_HVT U159 ( .A1(n66), .A2(n192), .Y(n68) );
  NAND2X0_HVT U160 ( .A1(n193), .A2(n68), .Y(n70) );
  INVX1_HVT U161 ( .A(n199), .Y(n65) );
  OAI21X1_HVT U162 ( .A1(n66), .A2(n201), .A3(n65), .Y(n67) );
  AOI21X1_HVT U163 ( .A1(n205), .A2(n68), .A3(n67), .Y(n69) );
  OAI21X1_HVT U164 ( .A1(n70), .A2(n207), .A3(n69), .Y(n73) );
  NAND2X0_HVT U165 ( .A1(n71), .A2(n196), .Y(n72) );
  XNOR2X1_HVT U166 ( .A1(n73), .A2(n72), .Y(sum[30]) );
  NOR2X0_HVT U167 ( .A1(n87), .A2(n192), .Y(n75) );
  NAND2X0_HVT U168 ( .A1(n193), .A2(n75), .Y(n77) );
  OAI21X1_HVT U169 ( .A1(n87), .A2(n201), .A3(n88), .Y(n74) );
  AOI21X1_HVT U170 ( .A1(n205), .A2(n75), .A3(n74), .Y(n76) );
  OAI21X1_HVT U171 ( .A1(n77), .A2(n207), .A3(n76), .Y(n82) );
  INVX1_HVT U172 ( .A(n78), .Y(n80) );
  NAND2X0_HVT U173 ( .A1(n80), .A2(n79), .Y(n81) );
  XNOR2X1_HVT U174 ( .A1(n82), .A2(n81), .Y(sum[29]) );
  INVX1_HVT U175 ( .A(n192), .Y(n84) );
  NAND2X0_HVT U176 ( .A1(n193), .A2(n84), .Y(n86) );
  INVX1_HVT U177 ( .A(n201), .Y(n83) );
  AOI21X1_HVT U178 ( .A1(n205), .A2(n84), .A3(n83), .Y(n85) );
  OAI21X1_HVT U179 ( .A1(n86), .A2(n207), .A3(n85), .Y(n91) );
  INVX1_HVT U180 ( .A(n87), .Y(n89) );
  NAND2X0_HVT U181 ( .A1(n89), .A2(n88), .Y(n90) );
  XNOR2X1_HVT U182 ( .A1(n91), .A2(n90), .Y(sum[28]) );
  INVX1_HVT U183 ( .A(n104), .Y(n92) );
  NOR2X0_HVT U184 ( .A1(n107), .A2(n92), .Y(n95) );
  NAND2X0_HVT U185 ( .A1(n193), .A2(n95), .Y(n97) );
  INVX1_HVT U186 ( .A(n103), .Y(n93) );
  OAI21X1_HVT U187 ( .A1(n107), .A2(n93), .A3(n108), .Y(n94) );
  AOI21X1_HVT U188 ( .A1(n205), .A2(n95), .A3(n94), .Y(n96) );
  OAI21X1_HVT U189 ( .A1(n97), .A2(n207), .A3(n96), .Y(n102) );
  INVX1_HVT U190 ( .A(n98), .Y(n100) );
  NAND2X0_HVT U191 ( .A1(n100), .A2(n99), .Y(n101) );
  XNOR2X1_HVT U192 ( .A1(n102), .A2(n101), .Y(sum[27]) );
  NAND2X0_HVT U193 ( .A1(n193), .A2(n104), .Y(n106) );
  AOI21X1_HVT U194 ( .A1(n205), .A2(n104), .A3(n103), .Y(n105) );
  OAI21X1_HVT U195 ( .A1(n106), .A2(n207), .A3(n105), .Y(n111) );
  INVX1_HVT U196 ( .A(n107), .Y(n109) );
  NAND2X0_HVT U197 ( .A1(n109), .A2(n108), .Y(n110) );
  XNOR2X1_HVT U198 ( .A1(n111), .A2(n110), .Y(sum[26]) );
  INVX1_HVT U199 ( .A(n112), .Y(n124) );
  NAND2X0_HVT U200 ( .A1(n193), .A2(n124), .Y(n115) );
  INVX1_HVT U201 ( .A(n123), .Y(n113) );
  AOI21X1_HVT U202 ( .A1(n205), .A2(n124), .A3(n113), .Y(n114) );
  OAI21X1_HVT U203 ( .A1(n115), .A2(n207), .A3(n114), .Y(n120) );
  INVX1_HVT U204 ( .A(n116), .Y(n118) );
  NAND2X0_HVT U205 ( .A1(n118), .A2(n117), .Y(n119) );
  XNOR2X1_HVT U206 ( .A1(n120), .A2(n119), .Y(sum[25]) );
  INVX1_HVT U207 ( .A(n193), .Y(n122) );
  INVX1_HVT U208 ( .A(n205), .Y(n121) );
  OAI21X1_HVT U209 ( .A1(n122), .A2(n207), .A3(n121), .Y(n126) );
  NAND2X0_HVT U210 ( .A1(n124), .A2(n123), .Y(n125) );
  XNOR2X1_HVT U211 ( .A1(n126), .A2(n125), .Y(sum[24]) );
  INVX1_HVT U212 ( .A(n159), .Y(n148) );
  INVX1_HVT U213 ( .A(n139), .Y(n127) );
  NOR2X0_HVT U214 ( .A1(n142), .A2(n127), .Y(n130) );
  NAND2X0_HVT U215 ( .A1(n148), .A2(n130), .Y(n132) );
  INVX1_HVT U216 ( .A(n158), .Y(n150) );
  INVX1_HVT U217 ( .A(n138), .Y(n128) );
  OAI21X1_HVT U218 ( .A1(n142), .A2(n128), .A3(n143), .Y(n129) );
  AOI21X1_HVT U219 ( .A1(n150), .A2(n130), .A3(n129), .Y(n131) );
  OAI21X1_HVT U220 ( .A1(n132), .A2(n207), .A3(n131), .Y(n137) );
  INVX1_HVT U221 ( .A(n133), .Y(n135) );
  NAND2X0_HVT U222 ( .A1(n135), .A2(n134), .Y(n136) );
  XNOR2X1_HVT U223 ( .A1(n137), .A2(n136), .Y(sum[23]) );
  NAND2X0_HVT U224 ( .A1(n148), .A2(n139), .Y(n141) );
  AOI21X1_HVT U225 ( .A1(n150), .A2(n139), .A3(n138), .Y(n140) );
  OAI21X1_HVT U226 ( .A1(n141), .A2(n207), .A3(n140), .Y(n146) );
  INVX1_HVT U227 ( .A(n142), .Y(n144) );
  NAND2X0_HVT U228 ( .A1(n144), .A2(n143), .Y(n145) );
  XNOR2X1_HVT U229 ( .A1(n146), .A2(n145), .Y(sum[22]) );
  INVX1_HVT U230 ( .A(n147), .Y(n161) );
  NAND2X0_HVT U231 ( .A1(n148), .A2(n161), .Y(n152) );
  INVX1_HVT U232 ( .A(n160), .Y(n149) );
  AOI21X1_HVT U233 ( .A1(n150), .A2(n161), .A3(n149), .Y(n151) );
  OAI21X1_HVT U234 ( .A1(n152), .A2(n207), .A3(n151), .Y(n157) );
  INVX1_HVT U235 ( .A(n153), .Y(n155) );
  NAND2X0_HVT U236 ( .A1(n155), .A2(n154), .Y(n156) );
  XNOR2X1_HVT U237 ( .A1(n157), .A2(n156), .Y(sum[21]) );
  OAI21X1_HVT U238 ( .A1(n159), .A2(n207), .A3(n158), .Y(n163) );
  NAND2X0_HVT U239 ( .A1(n161), .A2(n160), .Y(n162) );
  XNOR2X1_HVT U240 ( .A1(n163), .A2(n162), .Y(sum[20]) );
  INVX1_HVT U241 ( .A(n164), .Y(n178) );
  NAND2X0_HVT U242 ( .A1(n173), .A2(n178), .Y(n167) );
  INVX1_HVT U243 ( .A(n177), .Y(n165) );
  AOI21X1_HVT U244 ( .A1(n174), .A2(n178), .A3(n165), .Y(n166) );
  OAI21X1_HVT U245 ( .A1(n167), .A2(n207), .A3(n166), .Y(n172) );
  INVX1_HVT U246 ( .A(n168), .Y(n170) );
  NAND2X0_HVT U247 ( .A1(n170), .A2(n169), .Y(n171) );
  XNOR2X1_HVT U248 ( .A1(n172), .A2(n171), .Y(sum[19]) );
  INVX1_HVT U249 ( .A(n173), .Y(n176) );
  INVX1_HVT U250 ( .A(n174), .Y(n175) );
  OAI21X1_HVT U251 ( .A1(n176), .A2(n207), .A3(n175), .Y(n180) );
  NAND2X0_HVT U252 ( .A1(n178), .A2(n177), .Y(n179) );
  XNOR2X1_HVT U253 ( .A1(n180), .A2(n179), .Y(sum[18]) );
  OAI21X1_HVT U254 ( .A1(n186), .A2(n207), .A3(n187), .Y(n185) );
  INVX1_HVT U255 ( .A(n181), .Y(n183) );
  NAND2X0_HVT U256 ( .A1(n183), .A2(n182), .Y(n184) );
  XNOR2X1_HVT U257 ( .A1(n185), .A2(n184), .Y(sum[17]) );
  INVX1_HVT U258 ( .A(n186), .Y(n188) );
  NAND2X0_HVT U259 ( .A1(n188), .A2(n187), .Y(n189) );
  XOR2X1_HVT U260 ( .A1(n207), .A2(n189), .Y(sum[16]) );
  NOR2X0_HVT U261 ( .A1(n195), .A2(n190), .Y(n198) );
  NAND2X0_HVT U262 ( .A1(n191), .A2(n198), .Y(n202) );
  NOR2X0_HVT U263 ( .A1(n202), .A2(n192), .Y(n204) );
  NAND2X0_HVT U264 ( .A1(n193), .A2(n204), .Y(n208) );
  OAI21X1_HVT U265 ( .A1(n196), .A2(n195), .A3(n194), .Y(n197) );
  AOI21X1_HVT U266 ( .A1(n199), .A2(n198), .A3(n197), .Y(n200) );
  OAI21X1_HVT U267 ( .A1(n202), .A2(n201), .A3(n200), .Y(n203) );
  AOI21X1_HVT U268 ( .A1(n205), .A2(n204), .A3(n203), .Y(n206) );
  OAI21X1_HVT U269 ( .A1(n208), .A2(n207), .A3(n206), .Y(\intadd_0/n38 ) );
  INVX1_HVT U270 ( .A(n242), .Y(n231) );
  INVX1_HVT U271 ( .A(n222), .Y(n209) );
  NOR2X0_HVT U272 ( .A1(n225), .A2(n209), .Y(n213) );
  NAND2X0_HVT U273 ( .A1(n231), .A2(n213), .Y(n215) );
  INVX1_HVT U274 ( .A(n210), .Y(n273) );
  INVX1_HVT U275 ( .A(n241), .Y(n233) );
  INVX1_HVT U276 ( .A(n221), .Y(n211) );
  OAI21X1_HVT U277 ( .A1(n225), .A2(n211), .A3(n226), .Y(n212) );
  AOI21X1_HVT U278 ( .A1(n233), .A2(n213), .A3(n212), .Y(n214) );
  OAI21X1_HVT U279 ( .A1(n215), .A2(n273), .A3(n214), .Y(n220) );
  INVX1_HVT U280 ( .A(n216), .Y(n218) );
  NAND2X0_HVT U281 ( .A1(n218), .A2(n217), .Y(n219) );
  XNOR2X1_HVT U282 ( .A1(n220), .A2(n219), .Y(sum[15]) );
  NAND2X0_HVT U283 ( .A1(n231), .A2(n222), .Y(n224) );
  AOI21X1_HVT U284 ( .A1(n233), .A2(n222), .A3(n221), .Y(n223) );
  OAI21X1_HVT U285 ( .A1(n224), .A2(n273), .A3(n223), .Y(n229) );
  INVX1_HVT U286 ( .A(n225), .Y(n227) );
  NAND2X0_HVT U287 ( .A1(n227), .A2(n226), .Y(n228) );
  XNOR2X1_HVT U288 ( .A1(n229), .A2(n228), .Y(sum[14]) );
  INVX1_HVT U289 ( .A(n230), .Y(n244) );
  NAND2X0_HVT U290 ( .A1(n231), .A2(n244), .Y(n235) );
  INVX1_HVT U291 ( .A(n243), .Y(n232) );
  AOI21X1_HVT U292 ( .A1(n233), .A2(n244), .A3(n232), .Y(n234) );
  OAI21X1_HVT U293 ( .A1(n235), .A2(n273), .A3(n234), .Y(n240) );
  INVX1_HVT U294 ( .A(n236), .Y(n238) );
  NAND2X0_HVT U295 ( .A1(n238), .A2(n237), .Y(n239) );
  XNOR2X1_HVT U296 ( .A1(n240), .A2(n239), .Y(sum[13]) );
  OAI21X1_HVT U297 ( .A1(n242), .A2(n273), .A3(n241), .Y(n246) );
  NAND2X0_HVT U298 ( .A1(n244), .A2(n243), .Y(n245) );
  XNOR2X1_HVT U299 ( .A1(n246), .A2(n245), .Y(sum[12]) );
  INVX1_HVT U300 ( .A(n247), .Y(n261) );
  NAND2X0_HVT U301 ( .A1(n256), .A2(n261), .Y(n250) );
  INVX1_HVT U302 ( .A(n260), .Y(n248) );
  AOI21X1_HVT U303 ( .A1(n257), .A2(n261), .A3(n248), .Y(n249) );
  OAI21X1_HVT U304 ( .A1(n250), .A2(n273), .A3(n249), .Y(n255) );
  INVX1_HVT U305 ( .A(n251), .Y(n253) );
  NAND2X0_HVT U306 ( .A1(n253), .A2(n252), .Y(n254) );
  XNOR2X1_HVT U307 ( .A1(n255), .A2(n254), .Y(sum[11]) );
  INVX1_HVT U308 ( .A(n256), .Y(n259) );
  INVX1_HVT U309 ( .A(n257), .Y(n258) );
  OAI21X1_HVT U310 ( .A1(n259), .A2(n273), .A3(n258), .Y(n263) );
  NAND2X0_HVT U311 ( .A1(n261), .A2(n260), .Y(n262) );
  XNOR2X1_HVT U312 ( .A1(n263), .A2(n262), .Y(sum[10]) );
  OAI21X1_HVT U313 ( .A1(n269), .A2(n273), .A3(n270), .Y(n268) );
  INVX1_HVT U314 ( .A(n264), .Y(n266) );
  NAND2X0_HVT U315 ( .A1(n266), .A2(n265), .Y(n267) );
  XNOR2X1_HVT U316 ( .A1(n268), .A2(n267), .Y(sum[9]) );
  INVX1_HVT U317 ( .A(n269), .Y(n271) );
  NAND2X0_HVT U318 ( .A1(n271), .A2(n270), .Y(n272) );
  XOR2X1_HVT U319 ( .A1(n273), .A2(n272), .Y(sum[8]) );
  INVX1_HVT U320 ( .A(n274), .Y(n297) );
  AOI21X1_HVT U321 ( .A1(n297), .A2(n276), .A3(n275), .Y(n286) );
  OAI21X1_HVT U322 ( .A1(n282), .A2(n286), .A3(n283), .Y(n281) );
  INVX1_HVT U323 ( .A(n277), .Y(n279) );
  NAND2X0_HVT U324 ( .A1(n279), .A2(n278), .Y(n280) );
  XNOR2X1_HVT U325 ( .A1(n281), .A2(n280), .Y(sum[7]) );
  INVX1_HVT U326 ( .A(n282), .Y(n284) );
  NAND2X0_HVT U327 ( .A1(n284), .A2(n283), .Y(n285) );
  XOR2X1_HVT U328 ( .A1(n286), .A2(n285), .Y(sum[6]) );
  INVX1_HVT U329 ( .A(n287), .Y(n295) );
  INVX1_HVT U330 ( .A(n294), .Y(n288) );
  AOI21X1_HVT U331 ( .A1(n297), .A2(n295), .A3(n288), .Y(n293) );
  INVX1_HVT U332 ( .A(n289), .Y(n291) );
  NAND2X0_HVT U333 ( .A1(n291), .A2(n290), .Y(n292) );
  XOR2X1_HVT U334 ( .A1(n293), .A2(n292), .Y(sum[5]) );
  NAND2X0_HVT U335 ( .A1(n295), .A2(n294), .Y(n296) );
  XNOR2X1_HVT U336 ( .A1(n297), .A2(n296), .Y(sum[4]) );
  INVX1_HVT U337 ( .A(n298), .Y(n308) );
  OAI21X1_HVT U338 ( .A1(n304), .A2(n308), .A3(n305), .Y(n303) );
  INVX1_HVT U339 ( .A(n299), .Y(n301) );
  NAND2X0_HVT U340 ( .A1(n301), .A2(n300), .Y(n302) );
  XNOR2X1_HVT U341 ( .A1(n303), .A2(n302), .Y(sum[3]) );
  INVX1_HVT U342 ( .A(n304), .Y(n306) );
  NAND2X0_HVT U343 ( .A1(n306), .A2(n305), .Y(n307) );
  XOR2X1_HVT U344 ( .A1(n308), .A2(n307), .Y(sum[2]) );
  INVX1_HVT U345 ( .A(n309), .Y(n311) );
  NAND2X0_HVT U346 ( .A1(n311), .A2(n310), .Y(n313) );
  INVX1_HVT U347 ( .A(n314), .Y(n312) );
  XNOR2X1_HVT U348 ( .A1(n313), .A2(n312), .Y(sum[1]) );
  OA21X1_HVT U349 ( .A1(a[0]), .A2(b[0]), .A3(n314), .Y(sum[0]) );
endmodule
